`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/14/2019 12:11:14 PM
// Design Name: 
// Module Name: diff_io_mgr
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module dac_splitter #
  (
   parameter integer DATA_WIDTH = 14
   )
   (
	input clk,
	input rst,
	input dac_clk_i,
	input dac_wrt_i,
    input [DATA_WIDTH-1:0] 	din_a,
    input [DATA_WIDTH-1:0] 	din_b,
    output dac_clk_o,
    output dac_wrt_o,
    output dac_sel_o,
    output dac_rst_o,
	output [DATA_WIDTH-1:0] dout
    );

    ODDR ODDR_dac_clk ( .Q(dac_clk_o), .D1(1'b0), .D2(1'b1), .C(dac_clk_i),  .CE(1'b1), .R(rst), .S(1'b0) );
    ODDR ODDR_dac_wrt ( .Q(dac_wrt_o), .D1(1'b0), .D2(1'b1), .C(dac_wrt_i), .CE(1'b1), .R(rst), .S(1'b0) );
    ODDR ODDR_dac_sel ( .Q(dac_sel_o), .D1(1'b1), .D2(1'b0), .C(clk), .CE(1'b1), .R(rst), .S(1'b0) );
    ODDR ODDR_dac_rst ( .Q(dac_rst_o), .D1(rst), .D2(rst), .C(clk), .CE(1'b1), .R(1'b0), .S(1'b0) );
    
    ODDR ODDR_dac_0  ( .Q(dout[ 0]), .D1(din_b[ 0]), .D2(din_a[ 0]), .C(clk), .CE(1'b1), .R(rst), .S(1'b0) );
    ODDR ODDR_dac_1  ( .Q(dout[ 1]), .D1(din_b[ 1]), .D2(din_a[ 1]), .C(clk), .CE(1'b1), .R(rst), .S(1'b0) );
    ODDR ODDR_dac_2  ( .Q(dout[ 2]), .D1(din_b[ 2]), .D2(din_a[ 2]), .C(clk), .CE(1'b1), .R(rst), .S(1'b0) );
    ODDR ODDR_dac_3  ( .Q(dout[ 3]), .D1(din_b[ 3]), .D2(din_a[ 3]), .C(clk), .CE(1'b1), .R(rst), .S(1'b0) );
    ODDR ODDR_dac_4  ( .Q(dout[ 4]), .D1(din_b[ 4]), .D2(din_a[ 4]), .C(clk), .CE(1'b1), .R(rst), .S(1'b0) );
    ODDR ODDR_dac_5  ( .Q(dout[ 5]), .D1(din_b[ 5]), .D2(din_a[ 5]), .C(clk), .CE(1'b1), .R(rst), .S(1'b0) );
    ODDR ODDR_dac_6  ( .Q(dout[ 6]), .D1(din_b[ 6]), .D2(din_a[ 6]), .C(clk), .CE(1'b1), .R(rst), .S(1'b0) );
    ODDR ODDR_dac_7  ( .Q(dout[ 7]), .D1(din_b[ 7]), .D2(din_a[ 7]), .C(clk), .CE(1'b1), .R(rst), .S(1'b0) );
    ODDR ODDR_dac_8  ( .Q(dout[ 8]), .D1(din_b[ 8]), .D2(din_a[ 8]), .C(clk), .CE(1'b1), .R(rst), .S(1'b0) );
    ODDR ODDR_dac_9  ( .Q(dout[ 9]), .D1(din_b[ 9]), .D2(din_a[ 9]), .C(clk), .CE(1'b1), .R(rst), .S(1'b0) );
    ODDR ODDR_dac_10 ( .Q(dout[10]), .D1(din_b[10]), .D2(din_a[10]), .C(clk), .CE(1'b1), .R(rst), .S(1'b0) );
    ODDR ODDR_dac_11 ( .Q(dout[11]), .D1(din_b[11]), .D2(din_a[11]), .C(clk), .CE(1'b1), .R(rst), .S(1'b0) );
    ODDR ODDR_dac_12 ( .Q(dout[12]), .D1(din_b[12]), .D2(din_a[12]), .C(clk), .CE(1'b1), .R(rst), .S(1'b0) );
    ODDR ODDR_dac_13 ( .Q(dout[13]), .D1(din_b[13]), .D2(din_a[13]), .C(clk), .CE(1'b1), .R(rst), .S(1'b0) );
endmodule
